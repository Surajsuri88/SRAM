module tb;
reg clk;
reg rst;
reg[15:0]addr;
reg[15:0]wdata;
reg write;
reg valid;
wire[15:0]rdata;
wire ready;
wire error;
integer i;

Ram4Kb dut(clk,rst,addr,wdata,write,valid,rdata,error,ready);

//Clock Generation
initial begin
clk=0;
forever #5 clk=~clk;                           //10ns clock period
end

initial begin
rst=1; #15;
rst=0; 
end

//write operation
initial begin
#20;
for(i=0;i<=2047;i=i+1)begin

	addr=i;
	wdata=i+1;
	write=1;
	valid=1;
	#10;
end

rst=1;#10;

 //Read Operation
for(i=0;i<=2047;i=i+1)begin
	addr=i;
	write=0;
	valid=1;

	wait(ready==1)
	#10;
end
end

initial begin
$monitor(" addr=%d wdata=%d write=%d valid=%d rdata=%d ", addr,wdata,write,valid,rdata);
end
initial
#100000 $finish;

endmodule
